// Code your design here
module task_1(
  input [9:0]SW,
  output [9:0]LEDR
);
 assign LEDR = SW;
  
endmodule
  
